module lc3_output (
    input clk,
    input [7:0] data,
    input enable,
    output status

);

assign status = 1'b1;

endmodule